// Workaround BRAM implementation for fifo buffer
// 2020 <hackfin@section5.ch>

module bram_2psync_12_8_59fe624214af9b8daa183282288d5eb56b321f14 #(
	parameter DATA = 8,
	parameter ADDR = 12
) (

`include "bram.vh"


endmodule

module bram_2psync_6_8_59fe624214af9b8daa183282288d5eb56b321f14 #(
	parameter DATA = 8,
	parameter ADDR = 12
) (

`include "bram.vh"


endmodule
